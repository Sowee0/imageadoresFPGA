module CORR_SCORE(
	input				iCLK,
	input		[9:0] iPX_MEM,
	input		[9:0] iPX_REF,
	input		[9:0] iX,
	input		[9:0] iY,
	output	[9:0] oX,
	output 	[9:0]	oY
);
			


always @ (posedge iCLK) begin





end