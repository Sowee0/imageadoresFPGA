module SAVE_FRAME(

		input		iX,
		input		iY,
		input		iFrameCount,
		output 	oDone,
		output	oStopAck)
