module SAVE_FRAME(
				iRed,
				iGreen,
				iBlue,
				iSwitch,
				iX,
				iY,
				iCLK,
				oReady
				oStopcapture
				);
				

always @(posedge iCLK) begin

		if(iSwitch) begin
		
		
		
		end


end
				
