module IMG_SEARCH(

	input		[12:0]	iX,
	input 	[12:0] 	iY,
	output	[10:0] 	oVAL
	);
	
	parameter [3:0] halving = 4'd3; 
	
	reg 			decX;
	reg 			decY;
	reg 	[7:0] memPos;
	
	always @ (iX or iY) begin
	
	decX <= iX >> halving;
	decY <= iY >> halving;
	
	memPos =  decX + 12'd16 * decY;
	
	case (memPos)
		8d'0:		oVAL <= 10d'255;
		8d'1:		oVAL <= 10d'255;
		8d'2:		oVAL <= 10d'255;
		8d'3:		oVAL <= 10d'255;
		8d'4:		oVAL <= 10d'255;
		8d'5:		oVAL <= 10d'255;
		8d'6:		oVAL <= 10d'255;
		8d'7:		oVAL <= 10d'255;
		8d'8:		oVAL <= 10d'255;
		8d'9:		oVAL <= 10d'255;
		8d'10:	oVAL <= 10d'255;
		8d'11:	oVAL <= 10d'255;
		8d'12:	oVAL <= 10d'255;
		8d'13:	oVAL <= 10d'255;
		8d'14:	oVAL <= 10d'255;
		8d'15:	oVAL <= 10d'255;
		8d'16:	oVAL <= 10d'255;
		8d'17:	oVAL <= 10d'255;
		8d'18:	oVAL <= 10d'255;
		8d'19:	oVAL <= 10d'255;
		8d'20:	oVAL <= 10d'255;
		8d'21:	oVAL <= 10d'255;
		8d'22:	oVAL <= 10d'255;
		8d'23:	oVAL <= 10d'255;
		8d'24:	oVAL <= 10d'255;
		8d'25:	oVAL <= 10d'255;
		8d'26:	oVAL <= 10d'255;
		8d'27:	oVAL <= 10d'255;
		8d'28:	oVAL <= 10d'255;
		8d'29:	oVAL <= 10d'255;
		8d'30:	oVAL <= 10d'255;
		8d'31:	oVAL <= 10d'255;
		8d'32:	oVAL <= 10d'255;
		8d'33:	oVAL <= 10d'255;
		8d'34:	oVAL <= 10d'255;
		8d'35:	oVAL <= 10d'255;
		8d'36:	oVAL <= 10d'255;
		8d'37:	oVAL <= 10d'255;
		8d'38:	oVAL <= 10d'255;
		8d'39:	oVAL <= 10d'255;
		8d'40:	oVAL <= 10d'255;
		8d'41:	oVAL <= 10d'255;
		8d'42:	oVAL <= 10d'255;
		8d'43:	oVAL <= 10d'255;
		8d'44:	oVAL <= 10d'255;
		8d'45:	oVAL <= 10d'255;
		8d'46:	oVAL <= 10d'255;
		8d'47:	oVAL <= 10d'255;
		8d'48:	oVAL <= 10d'255;
		8d'49:	oVAL <= 10d'255;
		8d'50:	oVAL <= 10d'255;
		8d'51:	oVAL <= 10d'255;
		8d'52:	oVAL <= 10d'255;
		8d'53:	oVAL <= 10d'255;
		8d'54:	oVAL <= 10d'255;
		8d'55:	oVAL <= 10d'255;
		8d'56:	oVAL <= 10d'255;
		8d'57:	oVAL <= 10d'255;
		8d'58:	oVAL <= 10d'255;
		8d'59:	oVAL <= 10d'255;
		8d'60:	oVAL <= 10d'255;
		8d'61:	oVAL <= 10d'255;
		8d'62:	oVAL <= 10d'255;
		8d'63:	oVAL <= 10d'255;
		8d'64:	oVAL <= 10d'255;
		8d'65:	oVAL <= 10d'255;
		8d'66:	oVAL <= 10d'255;
		8d'67:	oVAL <= 10d'255;
		8d'68:	oVAL <= 10d'255;
		8d'69:	oVAL <= 10d'255;
		8d'70:	oVAL <= 10d'255;
		8d'71:	oVAL <= 10d'255;
		8d'72:	oVAL <= 10d'255;
		8d'73:	oVAL <= 10d'255;
		8d'74:	oVAL <= 10d'255;
		8d'75:	oVAL <= 10d'0;
		8d'76:	oVAL <= 10d'0;
		8d'77:	oVAL <= 10d'255;
		8d'78:	oVAL <= 10d'255;
		8d'79:	oVAL <= 10d'255;
		8d'80:	oVAL <= 10d'255;
		8d'81:	oVAL <= 10d'255;
		8d'82:	oVAL <= 10d'255;
		8d'83:	oVAL <= 10d'255;
		8d'84:	oVAL <= 10d'0;
		8d'85:	oVAL <= 10d'255;
		8d'86:	oVAL <= 10d'255;
		8d'87:	oVAL <= 10d'255;
		8d'88:	oVAL <= 10d'255;
		8d'89:	oVAL <= 10d'255;
		8d'90:	oVAL <= 10d'255;
		8d'91:	oVAL <= 10d'255;
		8d'92:	oVAL <= 10d'255;
		8d'93:	oVAL <= 10d'255;
		8d'94:	oVAL <= 10d'255;
		8d'95:	oVAL <= 10d'255;
		8d'96:	oVAL <= 10d'255;
		8d'97:	oVAL <= 10d'255;
		8d'98:	oVAL <= 10d'255;
		8d'99:	oVAL <= 10d'255;
		8d'100:	oVAL <= 10d'255;
		8d'101:	oVAL <= 10d'255;
		8d'102:	oVAL <= 10d'255;
		8d'103:	oVAL <= 10d'255;
		8d'104:	oVAL <= 10d'255;
		8d'105:	oVAL <= 10d'255;
		8d'106:	oVAL <= 10d'255;
		8d'107:	oVAL <= 10d'255;
		8d'108:	oVAL <= 10d'255;
		8d'109:	oVAL <= 10d'255;
		8d'110:	oVAL <= 10d'255;
		8d'111:	oVAL <= 10d'255;
		8d'112:	oVAL <= 10d'255;
		8d'113:	oVAL <= 10d'255;
		8d'114:	oVAL <= 10d'255;
		8d'115:	oVAL <= 10d'255;
		8d'116:	oVAL <= 10d'255;
		8d'117:	oVAL <= 10d'255;
		8d'118:	oVAL <= 10d'255;
		8d'119:	oVAL <= 10d'255;
		8d'120:	oVAL <= 10d'255;
		8d'121:	oVAL <= 10d'255;
		8d'122:	oVAL <= 10d'255;
		8d'123:	oVAL <= 10d'255;
		8d'124:	oVAL <= 10d'255;
		8d'125:	oVAL <= 10d'255;
		8d'126:	oVAL <= 10d'255;
		8d'127:	oVAL <= 10d'255;
		8d'128:	oVAL <= 10d'255;
		8d'129:	oVAL <= 10d'255;
		8d'130:	oVAL <= 10d'255;
		8d'131:	oVAL <= 10d'255;
		8d'132:	oVAL <= 10d'255;
		8d'133:	oVAL <= 10d'255;
		8d'134:	oVAL <= 10d'255;
		8d'135:	oVAL <= 10d'255;
		8d'136:	oVAL <= 10d'255;
		8d'137:	oVAL <= 10d'255;
		8d'138:	oVAL <= 10d'255;
		8d'139:	oVAL <= 10d'255;
		8d'140:	oVAL <= 10d'255;
		8d'141:	oVAL <= 10d'255;
		8d'142:	oVAL <= 10d'255;
		8d'143:	oVAL <= 10d'255;
		8d'144:	oVAL <= 10d'255;
		8d'145:	oVAL <= 10d'255;
		8d'146:	oVAL <= 10d'255;
		8d'147:	oVAL <= 10d'255;
		8d'148:	oVAL <= 10d'255;
		8d'149:	oVAL <= 10d'255;
		8d'150:	oVAL <= 10d'255;
		8d'151:	oVAL <= 10d'255;
		8d'152:	oVAL <= 10d'255;
		8d'153:	oVAL <= 10d'255;
		8d'154:	oVAL <= 10d'255;
		8d'155:	oVAL <= 10d'255;
		8d'156:	oVAL <= 10d'255;
		8d'157:	oVAL <= 10d'255;
		8d'158:	oVAL <= 10d'255;
		8d'159:	oVAL <= 10d'255;
		8d'160:	oVAL <= 10d'255;
		8d'161:	oVAL <= 10d'255;
		8d'162:	oVAL <= 10d'255;
		8d'163:	oVAL <= 10d'255;
		8d'164:	oVAL <= 10d'255;
		8d'165:	oVAL <= 10d'255;
		8d'166:	oVAL <= 10d'255;
		8d'167:	oVAL <= 10d'255;
		8d'168:	oVAL <= 10d'255;
		8d'169:	oVAL <= 10d'255;
		8d'170:	oVAL <= 10d'255;
		8d'171:	oVAL <= 10d'255;
		8d'172:	oVAL <= 10d'255;
		8d'173:	oVAL <= 10d'255;
		8d'174:	oVAL <= 10d'255;
		8d'175:	oVAL <= 10d'0;
		8d'176:	oVAL <= 10d'255;
		8d'177:	oVAL <= 10d'255;
		8d'178:	oVAL <= 10d'255;
		8d'179:	oVAL <= 10d'0;
		8d'180:	oVAL <= 10d'255;
		8d'181:	oVAL <= 10d'255;
		8d'182:	oVAL <= 10d'255;
		8d'183:	oVAL <= 10d'255;
		8d'184:	oVAL <= 10d'255;
		8d'185:	oVAL <= 10d'255;
		8d'186:	oVAL <= 10d'255;
		8d'187:	oVAL <= 10d'255;
		8d'188:	oVAL <= 10d'255;
		8d'189:	oVAL <= 10d'255;
		8d'190:	oVAL <= 10d'255;
		8d'191:	oVAL <= 10d'0;
		8d'192:	oVAL <= 10d'255;
		8d'193:	oVAL <= 10d'255;
		8d'194:	oVAL <= 10d'255;
		8d'195:	oVAL <= 10d'0;
		8d'196:	oVAL <= 10d'0;
		8d'197:	oVAL <= 10d'255;
		8d'198:	oVAL <= 10d'255;
		8d'199:	oVAL <= 10d'255;
		8d'200:	oVAL <= 10d'255;
		8d'201:	oVAL <= 10d'255;
		8d'202:	oVAL <= 10d'255;
		8d'203:	oVAL <= 10d'255;
		8d'204:	oVAL <= 10d'255;
		8d'205:	oVAL <= 10d'255;
		8d'206:	oVAL <= 10d'255;
		8d'207:	oVAL <= 10d'0;
		8d'208:	oVAL <= 10d'255;
		8d'209:	oVAL <= 10d'255;
		8d'210:	oVAL <= 10d'255;
		8d'211:	oVAL <= 10d'255;
		8d'212:	oVAL <= 10d'0;
		8d'213:	oVAL <= 10d'0;
		8d'214:	oVAL <= 10d'255;
		8d'215:	oVAL <= 10d'255;
		8d'216:	oVAL <= 10d'255;
		8d'217:	oVAL <= 10d'255;
		8d'218:	oVAL <= 10d'255;
		8d'219:	oVAL <= 10d'255;
		8d'220:	oVAL <= 10d'255;
		8d'221:	oVAL <= 10d'255;
		8d'222:	oVAL <= 10d'0;
		8d'223:	oVAL <= 10d'0;
		8d'224:	oVAL <= 10d'255;
		8d'225:	oVAL <= 10d'255;
		8d'226:	oVAL <= 10d'255;
		8d'227:	oVAL <= 10d'255;
		8d'228:	oVAL <= 10d'255;
		8d'229:	oVAL <= 10d'0;
		8d'230:	oVAL <= 10d'0;
		8d'231:	oVAL <= 10d'255;
		8d'232:	oVAL <= 10d'255;
		8d'233:	oVAL <= 10d'255;
		8d'234:	oVAL <= 10d'255;
		8d'235:	oVAL <= 10d'255;
		8d'236:	oVAL <= 10d'255;
		8d'237:	oVAL <= 10d'255;
		8d'238:	oVAL <= 10d'0;
		8d'239:	oVAL <= 10d'255;
		8d'240:	oVAL <= 10d'255;
		8d'241:	oVAL <= 10d'255;
		8d'242:	oVAL <= 10d'255;
		8d'243:	oVAL <= 10d'255;
		8d'244:	oVAL <= 10d'255;
		8d'245:	oVAL <= 10d'255;
		8d'246:	oVAL <= 10d'0;
		8d'247:	oVAL <= 10d'0;
		8d'248:	oVAL <= 10d'0;
		8d'249:	oVAL <= 10d'0;
		8d'250:	oVAL <= 10d'0;
		8d'251:	oVAL <= 10d'0;
		8d'252:	oVAL <= 10d'0;
		8d'253:	oVAL <= 10d'0;
		8d'254:	oVAL <= 10d'0;
		8d'255:	oVAL <= 10d'255;
		
		default: oVAL <= 10d'0;
		
		endcase

	end
	
	endmodule 