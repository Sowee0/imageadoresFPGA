// megafunction wizard: %Parallel Flash Loader%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altparallel_flash_loader 

// ============================================================
// File Name: tet.v
// Megafunction Name(s):
// 			altparallel_flash_loader
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
// ************************************************************

//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module tet (
	pfl_flash_access_granted,
	pfl_nreset,
	flash_addr,
	flash_data,
	flash_nce,
	flash_noe,
	flash_nwe,
	pfl_flash_access_request);

	input	  pfl_flash_access_granted;
	input	  pfl_nreset;
	output	[19:0]  flash_addr;
	inout	[7:0]  flash_data;
	output	  flash_nce;
	output	  flash_noe;
	output	  flash_nwe;
	output	  pfl_flash_access_request;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: DISABLE_CRC_CHECKBOX STRING "1"
// Retrieval info: PRIVATE: IDC_ENHANCED_FLASH_PROGRAMMING_COMBO STRING "Area"
// Retrieval info: PRIVATE: IDC_FIFO_SIZE_COMBO STRING "16"
// Retrieval info: PRIVATE: IDC_FLASH_DATA_WIDTH_COMBO STRING "8 bits"
// Retrieval info: PRIVATE: IDC_FLASH_DEVICE_COMBO STRING "CFI 8 Mbit"
// Retrieval info: PRIVATE: IDC_FLASH_NRESET_CHECKBOX STRING "0"
// Retrieval info: PRIVATE: IDC_FLASH_TYPE_COMBO STRING "CFI Parallel Flash"
// Retrieval info: PRIVATE: IDC_NUM_FLASH_COMBO STRING "1"
// Retrieval info: PRIVATE: IDC_OPERATING_MODES_COMBO STRING "Flash Programming"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: PRIVATE: TRISTATE_CHECKBOX STRING "0"
// Retrieval info: CONSTANT: ADDR_WIDTH NUMERIC "20"
// Retrieval info: CONSTANT: DISABLE_CRC_CHECKBOX NUMERIC "0"
// Retrieval info: CONSTANT: ENHANCED_FLASH_PROGRAMMING NUMERIC "0"
// Retrieval info: CONSTANT: FEATURES_CFG NUMERIC "0"
// Retrieval info: CONSTANT: FEATURES_PGM NUMERIC "1"
// Retrieval info: CONSTANT: FIFO_SIZE NUMERIC "16"
// Retrieval info: CONSTANT: FLASH_DATA_WIDTH NUMERIC "8"
// Retrieval info: CONSTANT: FLASH_NRESET_CHECKBOX NUMERIC "0"
// Retrieval info: CONSTANT: FLASH_TYPE STRING "CFI_FLASH"
// Retrieval info: CONSTANT: N_FLASH NUMERIC "1"
// Retrieval info: CONSTANT: TRISTATE_CHECKBOX NUMERIC "0"
// Retrieval info: USED_PORT: flash_addr 0 0 20 0 OUTPUT NODEFVAL "flash_addr[19..0]"
// Retrieval info: USED_PORT: flash_data 0 0 8 0 BIDIR NODEFVAL "flash_data[7..0]"
// Retrieval info: USED_PORT: flash_nce 0 0 0 0 OUTPUT NODEFVAL "flash_nce"
// Retrieval info: USED_PORT: flash_noe 0 0 0 0 OUTPUT NODEFVAL "flash_noe"
// Retrieval info: USED_PORT: flash_nwe 0 0 0 0 OUTPUT NODEFVAL "flash_nwe"
// Retrieval info: USED_PORT: pfl_flash_access_granted 0 0 0 0 INPUT NODEFVAL "pfl_flash_access_granted"
// Retrieval info: USED_PORT: pfl_flash_access_request 0 0 0 0 OUTPUT NODEFVAL "pfl_flash_access_request"
// Retrieval info: USED_PORT: pfl_nreset 0 0 0 0 INPUT NODEFVAL "pfl_nreset"
// Retrieval info: CONNECT: @pfl_flash_access_granted 0 0 0 0 pfl_flash_access_granted 0 0 0 0
// Retrieval info: CONNECT: @pfl_nreset 0 0 0 0 pfl_nreset 0 0 0 0
// Retrieval info: CONNECT: flash_addr 0 0 20 0 @flash_addr 0 0 20 0
// Retrieval info: CONNECT: flash_data 0 0 8 0 @flash_data 0 0 8 0
// Retrieval info: CONNECT: flash_nce 0 0 0 0 @flash_nce 0 0 0 0
// Retrieval info: CONNECT: flash_noe 0 0 0 0 @flash_noe 0 0 0 0
// Retrieval info: CONNECT: flash_nwe 0 0 0 0 @flash_nwe 0 0 0 0
// Retrieval info: CONNECT: pfl_flash_access_request 0 0 0 0 @pfl_flash_access_request 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL tet.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL tet.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL tet.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL tet.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL tet_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL tet_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
